
//------> /opt/catapult/Catapult_Synthesis_10.3d-815731/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /opt/catapult/Catapult_Synthesis_10.3d-815731/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /opt/catapult/Catapult_Synthesis_10.3d-815731/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.3d/815731 Production Release
//  HLS Date:       Wed Apr 24 14:54:19 PDT 2019
// 
//  Generated by:   student@SoC-courses
//  Generated date: Sat Mar 19 19:12:34 2022
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    determinant_core
// ------------------------------------------------------------------


module determinant_core (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, result_rsc_dat, result_rsc_triosy_lz
);
  input clk;
  input rst;
  input [152:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  output [16:0] result_rsc_dat;
  output result_rsc_triosy_lz;


  // Interconnect Declarations
  wire [152:0] input_rsci_idat;
  reg [16:0] result_rsci_idat;
  reg input_rsc_triosy_obj_ld;
  reg result_rsc_triosy_obj_ld;
  wire [1:0] determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp;
  wire [1:0] determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp;
  wire [1:0] determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_1_tmp;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_5_tmp;
  wire [2:0] input_mat_Matrix_for_1_for_acc_tmp;
  wire [4:0] nl_input_mat_Matrix_for_1_for_acc_tmp;
  wire and_dcpl;
  wire and_dcpl_1;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_12;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_17;
  wire and_dcpl_20;
  wire or_dcpl;
  wire and_dcpl_22;
  wire or_dcpl_4;
  wire nor_tmp;
  wire and_dcpl_26;
  wire and_dcpl_29;
  wire and_dcpl_32;
  wire and_dcpl_36;
  wire and_dcpl_48;
  wire and_dcpl_51;
  wire or_dcpl_10;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire and_dcpl_73;
  wire or_tmp_41;
  wire or_tmp_44;
  wire and_dcpl_89;
  wire and_dcpl_95;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire and_dcpl_109;
  wire or_dcpl_57;
  reg lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1;
  wire input_mat_Matrix_for_unequal_tmp_1;
  reg lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0;
  reg input_mat_Matrix_for_for_j_1_1_1_lpi_1;
  wire lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1;
  wire lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_or_m1c_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_3;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_28_cse_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_19_m1c_1;
  wire lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_2;
  reg [1:0] lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  wire lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1_1;
  wire lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0_1;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_or_47_ssc_1;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_26_ssc_1;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_27_ssc_1;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_25_ssc_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_25_ssc_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_44_ssc_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_or_3_tmp_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_or_1_psp_mx0;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_3;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_6_m1c_1;
  wire input_mat_Matrix_for_for_equal_tmp_2;
  wire input_mat_Matrix_for_for_equal_tmp_3;
  wire exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_4;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_14_ssc_1;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_and_15_ssc_1;
  wire exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_equal_tmp_2;
  wire input_mat_Matrix_for_i_1_1_lpi_1_dfm_1;
  wire input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1;
  wire input_mat_Matrix_for_for_or_m1c_1;
  wire lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_1_1;
  wire lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_0_1;
  reg input_mat_Matrix_for_asn_sft_lpi_1;
  wire lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1;
  wire input_mat_Matrix_for_for_and_ssc_1;
  wire input_mat_Matrix_for_for_and_6_ssc_1;
  wire lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_or_tmp_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_cse_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_cse_1;
  reg input_mat_Matrix_for_i_1_1_lpi_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_mx0;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_27_cse_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_2_tmp_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_tmp_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1;
  wire input_mat_Matrix_for_for_input_mat_Matrix_for_for_nor_3_cse_1;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_0;
  reg [1:0] lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_3;
  reg [1:0] lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_1_0;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_3;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_3;
  reg exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_3;
  reg [1:0] lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0;
  reg [1:0] lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_2;
  reg main_stage_0_3;
  reg [1:0] lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0;
  reg [1:0] lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  reg main_stage_0_2;
  reg [1:0] lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1;
  reg exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva;
  reg main_stage_0_4;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_3;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_2;
  reg exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_1;
  reg exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_1;
  reg sfi_exit_input_mat_Matrix_for_lpi_1;
  reg exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_4;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_0;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_1;
  reg main_stage_0_5;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_4;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_4;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_20_itm_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_11_itm_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_21_itm_1;
  wire [1:0] lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_dfm_4;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_41_itm_1;
  wire [1:0] lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_8_rgt;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_13_rgt;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_or_32_m1c;
  wire nor_11_cse;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_or_33_cse;
  wire and_124_cse;
  wire or_122_cse;
  wire determinant_helper_3_get_minor_ac_int_17_true_minor_data_or_1_cse;
  wire determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_3_cse;
  wire or_125_cse;
  wire and_123_cse;
  wire mux_15_cse;
  wire or_62_cse;
  wire or_22_cse;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_or_28_itm_1;
  reg [16:0] input_mat_data_1_2_lpi_1;
  reg [16:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_0_lpi_1;
  reg [16:0] input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1;
  reg [16:0] input_mat_data_2_0_lpi_1;
  wire [16:0] input_mat_data_2_1_lpi_1_mx0;
  wire and_128_tmp;
  wire or_127_tmp;
  wire mux_31_itm;
  wire and_dcpl_121;
  wire z_out_1;
  wire [30:0] z_out_3;
  wire [31:0] nl_z_out_3;
  reg [16:0] input_mat_data_1_1_lpi_1;
  reg [16:0] input_mat_data_1_0_lpi_1;
  reg [16:0] input_mat_data_0_2_lpi_1;
  reg [16:0] input_mat_data_0_1_lpi_1;
  reg [16:0] input_mat_data_2_1_lpi_1;
  reg [16:0] input_mat_data_0_0_lpi_1;
  reg [16:0] input_mat_data_2_2_lpi_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1;
  reg [16:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1;
  reg [16:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1;
  reg [29:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_31_2_lpi_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_lpi_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1;
  reg [16:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_dfm_6_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_dfm_1;
  reg [16:0] input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_4;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_2;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_3;
  reg [16:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_itm_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_acc_1_itm_1;
  wire [17:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_ac000000;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1;
  wire signed [34:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1;
  wire [17:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1;
  wire signed [33:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1;
  reg [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_acc_itm_1;
  reg [16:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_2_itm_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_40_itm_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_1;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_2;
  reg determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_3;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_3;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_1;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_2;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_3;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_4;
  reg determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_4;
  reg lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_1;
  wire result_rsci_idat_mx0c1;
  wire [16:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1;
  wire [17:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1;
  wire [16:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_mx0;
  wire [16:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_mx0;
  wire [16:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1_mx0;
  wire [16:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_2;
  wire [16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1_mx0;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_36_cse_mx0w0;
  wire [16:0] input_mat_data_2_2_lpi_1_mx0;
  wire [16:0] input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1_1;
  wire [16:0] input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_29_cse_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_and_30_cse_1;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_or_tmp_1;
  reg reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1_dfm_1_reg;
  reg reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg;
  wire determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_and_cse;
  wire input_mat_data_and_3_cse;
  wire nor_tmp_10;
  wire nor_tmp_15;
  wire not_tmp_119;
  wire or_tmp_77;
  wire nor_85_cse;
  wire nand_21_cse;
  wire nand_8_cse;
  wire nor_72_cse;
  wire and_182_cse;
  wire or_177_cse;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_itm_2;
  wire determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_itm_2;

  wire[0:0] mux_nl;
  wire[0:0] nor_43_nl;
  wire[0:0] nor_44_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] nor_41_nl;
  wire[0:0] nor_42_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nor_39_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] and_95_nl;
  wire[0:0] and_97_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] or_9_nl;
  wire[0:0] input_mat_Matrix_for_input_mat_Matrix_for_and_8_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_or_nl;
  wire[29:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_and_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_not_4_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_6_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_mux_4_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] or_130_nl;
  wire[0:0] and_187_nl;
  wire[0:0] or_129_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_9_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_or_1_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_12_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_2_nl;
  wire[1:0] determinant_helper_3_do_determinant_ac_int_17_true_for_and_28_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_nor_1_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] and_120_nl;
  wire[0:0] and_121_nl;
  wire[0:0] or_17_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] or_15_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_mux_4_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_or_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_nor_1_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] nand_20_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] nor_79_nl;
  wire[0:0] or_178_nl;
  wire[0:0] input_mat_Matrix_for_not_17_nl;
  wire[0:0] input_mat_Matrix_for_for_input_mat_Matrix_for_for_mux_22_nl;
  wire[16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_nl;
  wire signed [33:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_nl;
  wire[16:0] determinant_helper_2_do_determinant_ac_int_17_true_for_mux_6_nl;
  wire[16:0] determinant_helper_2_do_determinant_ac_int_17_true_for_mux_7_nl;
  wire[16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_nl;
  wire signed [33:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_nl;
  wire[0:0] and_100_nl;
  wire[0:0] and_101_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] nor_73_nl;
  wire[0:0] nor_74_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_52_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_or_26_nl;
  wire[0:0] mux_51_nl;
  wire[0:0] or_153_nl;
  wire[0:0] mux_50_nl;
  wire[0:0] mux_49_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] and_184_nl;
  wire[0:0] or_150_nl;
  wire[16:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_1_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_45_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_or_25_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_48_nl;
  wire[0:0] mux_58_nl;
  wire[0:0] nand_13_nl;
  wire[0:0] mux_57_nl;
  wire[0:0] mux_56_nl;
  wire[0:0] or_161_nl;
  wire[0:0] mux_55_nl;
  wire[0:0] mux_54_nl;
  wire[0:0] or_160_nl;
  wire[0:0] mux_53_nl;
  wire[0:0] or_159_nl;
  wire[0:0] or_158_nl;
  wire[0:0] mux_52_nl;
  wire[0:0] and_183_nl;
  wire[0:0] or_155_nl;
  wire[0:0] or_154_nl;
  wire[16:0] mux1h_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_33_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_56_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_and_57_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_and_35_nl;
  wire[0:0] not_235_nl;
  wire[0:0] mux_65_nl;
  wire[0:0] or_179_nl;
  wire[0:0] or_180_nl;
  wire[0:0] mux_64_nl;
  wire[0:0] mux_63_nl;
  wire[0:0] nor_82_nl;
  wire[0:0] mux_62_nl;
  wire[0:0] nor_83_nl;
  wire[0:0] or_169_nl;
  wire[0:0] mux_61_nl;
  wire[0:0] mux_60_nl;
  wire[0:0] or_168_nl;
  wire[0:0] or_167_nl;
  wire[0:0] mux_59_nl;
  wire[0:0] nand_23_nl;
  wire[0:0] or_166_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] or_73_nl;
  wire[0:0] or_71_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] nor_15_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] nor_16_nl;
  wire[16:0] determinant_helper_3_do_determinant_ac_int_17_true_for_2_acc_1_nl;
  wire[17:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_2_acc_1_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_or_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_and_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_determinant_and_1_nl;
  wire[2:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_nl;
  wire[4:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_nl;
  wire[31:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_nl;
  wire[32:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_nl;
  wire[2:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_nl;
  wire[4:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_and_29_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_and_30_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_or_30_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_2_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_for_not_30_nl;
  wire[0:0] determinant_helper_3_do_determinant_ac_int_17_true_for_mux_5_nl;
  wire[0:0] input_mat_Matrix_for_for_mux_20_nl;
  wire[0:0] input_mat_Matrix_for_for_input_mat_Matrix_for_nor_nl;
  wire[2:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_nl;
  wire[4:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_nl;
  wire[2:0] determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_nl;
  wire[4:0] nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_nl;
  wire[0:0] determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_2_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] or_47_nl;
  wire[0:0] or_46_nl;
  wire[16:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_8_nl;
  wire[16:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_4_nl;
  wire[0:0] nor_48_nl;
  wire[0:0] and_134_nl;
  wire[16:0] determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_6_nl;
  wire[0:0] asn_input_mat_data_2_1_lpi_1_nand_nl;
  wire[0:0] asn_input_mat_data_2_2_lpi_1_nand_nl;
  wire[0:0] or_108_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] nor_25_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] or_31_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] or_29_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] nor_29_nl;
  wire[0:0] nor_86_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] nor_19_nl;
  wire[30:0] determinant_helper_3_do_determinant_ac_int_17_true_for_mux_15_nl;
  wire[0:0] input_mat_Matrix_for_for_mux_25_nl;
  wire[0:0] input_mat_Matrix_for_for_input_mat_Matrix_for_for_or_6_nl;
  wire[0:0] input_mat_Matrix_for_for_mux_26_nl;

  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd153)) input_rsci (
      .dat(input_rsc_dat),
      .idat(input_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd2),
  .width(32'sd17)) result_rsci (
      .idat(result_rsci_idat),
      .dat(result_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_rsc_triosy_obj (
      .ld(input_rsc_triosy_obj_ld),
      .lz(input_rsc_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) result_rsc_triosy_obj (
      .ld(result_rsc_triosy_obj_ld),
      .lz(result_rsc_triosy_lz)
    );
  assign nor_11_cse = ~((determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp!=2'b00));
  assign nor_85_cse = ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_and_cse = or_dcpl_4
      & (~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | or_dcpl));
  assign nand_21_cse = ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
      & (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_33_cse = (mux_15_cse
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0))
      | and_dcpl_109;
  assign nor_72_cse = ~(and_124_cse | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign or_177_cse = nor_72_cse | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva;
  assign nand_8_cse = ~(determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1);
  assign and_182_cse = determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_32_m1c = determinant_helper_3_get_minor_ac_int_17_true_for_and_36_cse_mx0w0
      | ((~(determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1 | (~
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2)))
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1);
  assign or_125_cse = (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp!=2'b00);
  assign and_128_tmp = (~((~((~((~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2)
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1))
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1)) & determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_3))
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign and_124_cse = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign or_62_cse = (input_mat_Matrix_for_1_for_acc_tmp[2:1]!=2'b00);
  assign or_122_cse = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 | input_mat_Matrix_for_for_j_1_1_1_lpi_1;
  assign or_73_nl = (~(lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 | input_mat_Matrix_for_i_1_1_lpi_1))
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1;
  assign mux_33_nl = MUX_s_1_2_2((or_73_nl), or_tmp_41, lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0);
  assign or_71_nl = and_123_cse | (~ input_mat_Matrix_for_i_1_1_lpi_1) | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1;
  assign mux_34_nl = MUX_s_1_2_2((mux_33_nl), (or_71_nl), input_mat_Matrix_for_asn_sft_lpi_1);
  assign mux_35_nl = MUX_s_1_2_2((~ mux_31_itm), (mux_34_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign input_mat_data_and_3_cse = (~((mux_35_nl) | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva))
      & (~(or_dcpl_57 | (~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
      & sfi_exit_input_mat_Matrix_for_lpi_1))));
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1
      = determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1 +
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1 = nl_determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1[16:0];
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_2_acc_1_nl = determinant_helper_3_do_determinant_ac_int_17_true_determinant_lpi_1
      + determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_2_acc_1_nl = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_2_acc_1_nl[16:0];
  assign determinant_helper_3_do_determinant_ac_int_17_true_determinant_or_nl = (~
      main_stage_0_5) | determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_4;
  assign determinant_helper_3_do_determinant_ac_int_17_true_determinant_and_nl =
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_4 & main_stage_0_5;
  assign determinant_helper_3_do_determinant_ac_int_17_true_determinant_and_1_nl
      = determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_4 & main_stage_0_5;
  assign determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_mx0
      = MUX1HOT_v_17_3_2(determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1,
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_dfm_1,
      (determinant_helper_3_do_determinant_ac_int_17_true_for_2_acc_1_nl), {(determinant_helper_3_do_determinant_ac_int_17_true_determinant_or_nl)
      , (determinant_helper_3_do_determinant_ac_int_17_true_determinant_and_nl) ,
      (determinant_helper_3_do_determinant_ac_int_17_true_determinant_and_1_nl)});
  assign lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1
      = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
      & determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_2;
  assign lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1
      = MUX_v_2_2_2(2'b00, lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0,
      determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_2);
  assign exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2 = input_mat_Matrix_for_i_1_1_lpi_1_dfm_1
      & input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1 & input_mat_Matrix_for_for_or_m1c_1;
  assign lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
      & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1
      = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
      & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1 = input_mat_Matrix_for_for_j_1_1_1_lpi_1
      & input_mat_Matrix_for_unequal_tmp_1;
  assign lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1 = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1
      & input_mat_Matrix_for_unequal_tmp_1;
  assign lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1 = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0
      & input_mat_Matrix_for_unequal_tmp_1;
  assign input_mat_Matrix_for_unequal_tmp_1 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1
      & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1==2'b00);
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_nl
      = ({1'b1 , (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      , 1'b1}) + conv_u2s_2_3({determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1
      , 1'b0}) + 3'b001;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_nl[2:0];
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2
      = readslicef_3_1_2((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_nl));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1
      = determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1 & determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_2;
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_nl
      = ({determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_31_2_lpi_1
      , determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1 ,
      1'b1}) + 32'b11111111111111111111111111111101;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_nl[31:0];
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31
      = readslicef_32_1_31((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_nl));
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_nl
      = ({1'b1 , (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      , 1'b1}) + conv_u2s_2_3({determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1
      , 1'b0}) + 3'b001;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_nl[2:0];
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2
      = readslicef_3_1_2((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_nl));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_13_rgt = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_2 = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1!=2'b00);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_29_nl = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1)
      & determinant_helper_3_do_determinant_ac_int_17_true_for_and_25_ssc_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_30_nl = determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_and_25_ssc_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_1_tmp
      = MUX1HOT_v_2_4_2(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0,
      2'b01, 2'b10, lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1,
      {determinant_helper_3_do_determinant_ac_int_17_true_for_or_47_ssc_1 , (determinant_helper_3_do_determinant_ac_int_17_true_for_and_29_nl)
      , (determinant_helper_3_do_determinant_ac_int_17_true_for_and_30_nl) , determinant_helper_3_do_determinant_ac_int_17_true_for_and_26_ssc_1});
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp = MUX_v_2_2_2((signext_2_1(~
      exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2)), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_dfm_4,
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2);
  assign exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_4
      = determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3 & determinant_helper_3_get_minor_ac_int_17_true_for_or_m1c_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_3;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_m1c_1 = ((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1==2'b01))
      | (~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1!=2'b00)));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_3 = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_dfm_4!=2'b00);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_30_nl = ((~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3)
      & determinant_helper_3_get_minor_ac_int_17_true_for_or_m1c_1) | determinant_helper_3_get_minor_ac_int_17_true_for_and_28_cse_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_2_nl
      = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1==2'b11);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp = MUX1HOT_v_2_3_2(2'b01,
      2'b10, lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1,
      {(determinant_helper_3_get_minor_ac_int_17_true_for_or_30_nl) , determinant_helper_3_get_minor_ac_int_17_true_for_and_27_cse_1
      , (determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_2_nl)});
  assign determinant_helper_3_get_minor_ac_int_17_true_for_not_30_nl = ~ determinant_helper_3_get_minor_ac_int_17_true_for_equal_tmp_2;
  assign lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_dfm_4
      = MUX_v_2_2_2(2'b00, determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp,
      (determinant_helper_3_get_minor_ac_int_17_true_for_not_30_nl));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_28_cse_1 = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_19_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_27_cse_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_19_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_equal_tmp_2 = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1==2'b10);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_19_m1c_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_mux_5_nl = MUX_s_1_2_2((~
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_4), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1,
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_3);
  assign lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1_1
      = ((determinant_helper_3_do_determinant_ac_int_17_true_for_mux_5_nl) & (~ determinant_helper_3_do_determinant_ac_int_17_true_for_and_14_ssc_1))
      | determinant_helper_3_do_determinant_ac_int_17_true_for_and_15_ssc_1;
  assign lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0_1
      = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1
      & (~(determinant_helper_3_do_determinant_ac_int_17_true_for_and_15_ssc_1 |
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2))) | determinant_helper_3_do_determinant_ac_int_17_true_for_and_14_ssc_1;
  assign input_mat_Matrix_for_for_input_mat_Matrix_for_nor_nl = ~((~ sfi_exit_input_mat_Matrix_for_lpi_1)
      | input_mat_Matrix_for_asn_sft_lpi_1);
  assign input_mat_Matrix_for_for_mux_20_nl = MUX_s_1_2_2((input_mat_Matrix_for_for_input_mat_Matrix_for_nor_nl),
      lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1, input_mat_Matrix_for_for_equal_tmp_3);
  assign lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_1_1 = ((input_mat_Matrix_for_for_mux_20_nl)
      & (~ input_mat_Matrix_for_for_and_ssc_1)) | input_mat_Matrix_for_for_and_6_ssc_1;
  assign lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_0_1 = (lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1
      & (~(input_mat_Matrix_for_for_and_6_ssc_1 | input_mat_Matrix_for_for_equal_tmp_2)))
      | input_mat_Matrix_for_for_and_ssc_1;
  assign input_mat_Matrix_for_i_1_1_lpi_1_dfm_1 = input_mat_Matrix_for_i_1_1_lpi_1
      & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign input_mat_Matrix_for_for_equal_tmp_2 = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1
      & (~ lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1);
  assign input_mat_Matrix_for_for_equal_tmp_3 = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1
      & lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1 = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1))
      | (~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1));
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_3 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_or_47_ssc_1 = (~
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2) | determinant_helper_3_get_minor_ac_int_17_true_for_or_1_psp_mx0;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_26_ssc_1 = ((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1) | (determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1
      & (~ determinant_helper_3_get_minor_ac_int_17_true_for_or_1_psp_mx0)) | determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1)
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_27_ssc_1 = determinant_helper_3_get_minor_ac_int_17_true_for_and_19_m1c_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_25_ssc_1 = determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_25_ssc_1 = (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31)
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_44_ssc_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_or_3_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1 = ~(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_itm_2
      & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_or_3_tmp_1 = ~(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_itm_2
      & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1 = ~(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_cse_1
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_cse_1
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4 | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_1_psp_mx0 = MUX_s_1_2_2((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]),
      determinant_helper_3_get_minor_ac_int_17_true_for_and_40_itm_1, or_dcpl_41);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_or_tmp_1
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_nl
      = ({1'b1 , (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      , 1'b1}) + conv_u2s_2_3({determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1
      , 1'b1}) + 3'b001;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_nl[2:0];
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_itm_2
      = readslicef_3_1_2((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_nl));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4 = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1[1])
      & (~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1[0])));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5 = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1==2'b11)
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_8_rgt = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_or_tmp_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_cse_1
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_cse_1;
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_nl
      = ({1'b1 , (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      , 1'b1}) + conv_u2s_2_3({determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1
      , 1'b1}) + 3'b001;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_nl[2:0];
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_itm_2
      = readslicef_3_1_2((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_nl));
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_5_tmp = (~ determinant_helper_3_get_minor_ac_int_17_true_for_equal_tmp_2)
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_6_m1c_1 = determinant_helper_3_get_minor_ac_int_17_true_for_equal_tmp_2
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign input_mat_Matrix_for_for_input_mat_Matrix_for_for_nor_3_cse_1 = ~(input_mat_Matrix_for_for_equal_tmp_2
      | input_mat_Matrix_for_for_equal_tmp_3);
  assign input_mat_Matrix_for_for_or_m1c_1 = (lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1
      & (~ lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1)) | (~(lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_1_1
      | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_0_1));
  assign input_mat_Matrix_for_for_and_ssc_1 = (~ input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1)
      & input_mat_Matrix_for_for_or_m1c_1;
  assign input_mat_Matrix_for_for_and_6_ssc_1 = input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1
      & input_mat_Matrix_for_for_or_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_cse_1
      = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1[0])
      & (~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1[1])));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_cse_1
      = ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1!=2'b00));
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_14_ssc_1 = (~
      exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2) & determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1;
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_15_ssc_1 = exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2
      & determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_minor_data_or_1_cse = (~ main_stage_0_2)
      | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_3_cse = determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1
      & main_stage_0_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_2_nl = determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1
      & main_stage_0_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_mx0 =
      MUX1HOT_v_17_3_2(determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1,
      ({{16{reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg}},
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg}),
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_dfm_6_1,
      {determinant_helper_3_get_minor_ac_int_17_true_minor_data_or_1_cse , (determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_2_nl)
      , determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_3_cse});
  assign or_127_tmp = (determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_or_28_itm_1 & determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_3_cse)
      | determinant_helper_3_get_minor_ac_int_17_true_minor_data_or_1_cse;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_4_nl
      = MUX1HOT_v_17_3_2(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1,
      input_mat_data_2_1_lpi_1, input_mat_data_2_2_lpi_1, {determinant_helper_3_get_minor_ac_int_17_true_for_and_40_itm_1
      , determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1_1 , determinant_helper_3_get_minor_ac_int_17_true_for_and_41_itm_1});
  assign determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_8_nl
      = MUX_v_17_2_2(17'b00000000000000000, (determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_4_nl),
      determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1);
  assign nor_48_nl = ~(determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_3_cse
      | or_127_tmp);
  assign and_134_nl = determinant_helper_3_get_minor_ac_int_17_true_minor_data_and_3_cse
      & (~ or_127_tmp);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1_mx0
      = MUX1HOT_v_17_3_2(({{16{reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1_dfm_1_reg}},
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1_dfm_1_reg}),
      (determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_8_nl),
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1, {(nor_48_nl)
      , (and_134_nl) , or_127_tmp});
  assign determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_6_nl
      = MUX_v_17_2_2(17'b00000000000000000, determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_2_itm_1,
      determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1);
  assign determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_2 = MUX_v_17_2_2(({{16{reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg}},
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg}),
      (determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_and_6_nl),
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1_mx0
      = MUX_v_17_2_2(input_mat_data_1_0_lpi_1, input_mat_data_1_2_lpi_1, z_out_3[0]);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_36_cse_mx0w0 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_2_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1;
  assign asn_input_mat_data_2_1_lpi_1_nand_nl = ~(main_stage_0_2 & determinant_helper_3_do_determinant_ac_int_17_true_for_and_11_itm_1);
  assign input_mat_data_2_1_lpi_1_mx0 = MUX_v_17_2_2(input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1,
      input_mat_data_2_1_lpi_1, asn_input_mat_data_2_1_lpi_1_nand_nl);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1 = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_or_3_tmp_1)
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1;
  assign asn_input_mat_data_2_2_lpi_1_nand_nl = ~(main_stage_0_2 & determinant_helper_3_do_determinant_ac_int_17_true_for_and_21_itm_1);
  assign input_mat_data_2_2_lpi_1_mx0 = MUX_v_17_2_2(input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1,
      input_mat_data_2_2_lpi_1, asn_input_mat_data_2_2_lpi_1_nand_nl);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3;
  assign or_108_nl = or_dcpl | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_mx0 =
      MUX_s_1_2_2(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_1,
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp, or_108_nl);
  assign input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1_1
      = MUX_v_17_5_2((input_rsci_idat[16:0]), (input_rsci_idat[50:34]), (input_rsci_idat[84:68]),
      (input_rsci_idat[118:102]), (input_rsci_idat[152:136]), input_mat_Matrix_for_1_for_acc_tmp);
  assign input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1_1
      = MUX_v_17_4_2x1x2((input_rsci_idat[33:17]), (input_rsci_idat[135:119]), {{1{input_mat_Matrix_for_i_1_1_lpi_1_dfm_1}},
      input_mat_Matrix_for_i_1_1_lpi_1_dfm_1});
  assign nl_input_mat_Matrix_for_1_for_acc_tmp = conv_u2u_2_3({input_mat_Matrix_for_i_1_1_lpi_1_dfm_1
      , 1'b0}) + conv_u2u_1_3(input_mat_Matrix_for_i_1_1_lpi_1_dfm_1) + conv_u2u_1_3(input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1);
  assign input_mat_Matrix_for_1_for_acc_tmp = nl_input_mat_Matrix_for_1_for_acc_tmp[2:0];
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_2_tmp_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_29_cse_1 = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_tmp_1)
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_30_cse_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_or_tmp_1 = determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_tmp_1 = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1)
      & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31;
  assign and_dcpl = main_stage_0_4 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_1;
  assign and_dcpl_1 = and_dcpl & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_0);
  assign and_dcpl_9 = main_stage_0_3 & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0);
  assign and_dcpl_10 = and_dcpl_9 & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2[1]))
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1;
  assign and_dcpl_12 = and_dcpl_9 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1;
  assign and_dcpl_14 = main_stage_0_2 & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0);
  assign and_dcpl_15 = and_dcpl_14 & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[1]))
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1;
  assign and_dcpl_17 = and_dcpl_14 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1;
  assign and_dcpl_20 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      & nor_85_cse;
  assign or_dcpl = exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign and_dcpl_22 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign and_123_cse = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 & lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0;
  assign or_dcpl_4 = (~(and_123_cse | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1))
      | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva | (~
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign nor_tmp = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 & lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign or_22_cse = nor_11_cse | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1) | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00);
  assign nor_27_nl = ~((~ determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_2)
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2!=2'b10));
  assign nor_28_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2[1])
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0[1])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0[0]));
  assign mux_13_nl = MUX_s_1_2_2((nor_27_nl), (nor_28_nl), determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_2);
  assign and_dcpl_26 = (mux_13_nl) & and_dcpl_12;
  assign nor_25_nl = ~((~ determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_1)
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1!=2'b10));
  assign nor_26_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[1])
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0[1])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0[0]));
  assign mux_14_nl = MUX_s_1_2_2((nor_25_nl), (nor_26_nl), determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_1);
  assign and_dcpl_29 = (mux_14_nl) & and_dcpl_17;
  assign or_31_nl = (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]));
  assign mux_15_cse = MUX_s_1_2_2((or_31_nl), (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]),
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]);
  assign or_29_nl = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]));
  assign mux_16_nl = MUX_s_1_2_2(mux_15_cse, (or_29_nl), determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1);
  assign and_dcpl_32 = (~ (mux_16_nl)) & and_dcpl_22;
  assign and_dcpl_36 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
      & (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign and_dcpl_48 = ~(nor_72_cse | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign and_dcpl_51 = determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_and_5_tmp;
  assign or_dcpl_10 = (determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp!=2'b10);
  assign and_dcpl_68 = ~(exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign and_dcpl_69 = and_dcpl_68 & input_mat_Matrix_for_i_1_1_lpi_1;
  assign nor_29_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1));
  assign mux_11_nl = MUX_s_1_2_2((nor_29_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1,
      or_22_cse);
  assign nor_86_nl = ~((~ input_mat_Matrix_for_for_j_1_1_1_lpi_1) | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1
      | (~ input_mat_Matrix_for_i_1_1_lpi_1) | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign mux_12_nl = MUX_s_1_2_2((mux_11_nl), (nor_86_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign and_dcpl_73 = (mux_12_nl) & or_dcpl_10 & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign or_tmp_41 = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 | (~ input_mat_Matrix_for_i_1_1_lpi_1)
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1;
  assign or_tmp_44 = input_mat_Matrix_for_i_1_1_lpi_1 | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1;
  assign nor_19_nl = ~((~ input_mat_Matrix_for_i_1_1_lpi_1) | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign mux_30_nl = MUX_s_1_2_2(or_tmp_44, (nor_19_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign mux_31_itm = MUX_s_1_2_2((mux_30_nl), or_tmp_44, or_22_cse);
  assign and_dcpl_89 = main_stage_0_5 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_1
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_0);
  assign and_dcpl_95 = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
      & (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign or_dcpl_41 = or_dcpl | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign or_dcpl_42 = ~(main_stage_0_2 & determinant_helper_3_do_determinant_ac_int_17_true_for_and_20_itm_1);
  assign and_dcpl_109 = and_dcpl_95 & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0==2'b00)
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1 &
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
      & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]))
      & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign or_dcpl_57 = (~ lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1) | input_mat_Matrix_for_asn_sft_lpi_1;
  assign result_rsci_idat_mx0c1 = and_dcpl_89 & exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_4
      & (~ determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_4);
  assign and_dcpl_121 = lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign nor_tmp_10 = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2
      & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_itm_2;
  assign nor_tmp_15 = determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1;
  assign not_tmp_119 = determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1
      & nor_tmp_15;
  assign or_tmp_77 = (~ main_stage_0_2) | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  always @(posedge clk) begin
    if ( rst ) begin
      result_rsc_triosy_obj_ld <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_1
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_0
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_1
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_0
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0
          <= 1'b0;
      input_rsc_triosy_obj_ld <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
          <= 1'b0;
      exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva <= 1'b1;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
          <= 1'b0;
      main_stage_0_2 <= 1'b0;
      main_stage_0_3 <= 1'b0;
      main_stage_0_4 <= 1'b0;
      main_stage_0_5 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_4 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_4 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_4 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_4 <= 1'b0;
      input_mat_Matrix_for_i_1_1_lpi_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_3 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_3 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_3 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_3 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_2 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_2 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_2 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_2 <= 1'b0;
      determinant_helper_3_get_minor_ac_int_17_true_for_or_28_itm_1 <= 1'b0;
      determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_21_itm_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_20_itm_1 <= 1'b0;
    end
    else begin
      result_rsc_triosy_obj_ld <= main_stage_0_5 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_1
          & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_0)
          & exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_4;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_1
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_1;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_4_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_1
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_0_1;
      input_rsc_triosy_obj_ld <= ~((~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1)
          | (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]))
          | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
          | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
          | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
          | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
          | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva
          | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
          | nor_11_cse | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1_1;
      exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva <= ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1_1
          | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0_1);
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0_1;
      main_stage_0_2 <= 1'b1;
      main_stage_0_3 <= main_stage_0_2;
      main_stage_0_4 <= main_stage_0_3;
      main_stage_0_5 <= main_stage_0_4;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_4 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_3;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_4 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_3;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_4 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_3;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_4 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_3;
      input_mat_Matrix_for_i_1_1_lpi_1 <= MUX_s_1_2_2(input_mat_Matrix_for_i_1_1_lpi_1_dfm_1,
          (input_mat_Matrix_for_for_input_mat_Matrix_for_for_mux_22_nl), or_dcpl);
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_3 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_3 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_3 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_3 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_2 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_2 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_2 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_2 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
      determinant_helper_3_get_minor_ac_int_17_true_for_or_28_itm_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_for_1_or_tmp_1
          | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1 | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
          | ((~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_2_tmp_1)
          & determinant_helper_3_get_minor_ac_int_17_true_for_and_10_m1c_1) | determinant_helper_3_get_minor_ac_int_17_true_for_and_27_cse_1
          | (determinant_helper_3_get_minor_ac_int_17_true_for_for_or_3_tmp_1 & determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1);
      determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_and_54_itm_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1 <= determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_1 <= (~ determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1)
          & determinant_helper_3_do_determinant_ac_int_17_true_for_and_6_m1c_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_1 <= determinant_helper_3_do_determinant_ac_int_17_true_for_and_5_tmp
          | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_3 |
          (determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1 &
          determinant_helper_3_do_determinant_ac_int_17_true_for_and_6_m1c_1);
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_mx0
          & (~ determinant_helper_3_get_minor_ac_int_17_true_for_or_1_psp_mx0) &
          determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_21_itm_1 <= (input_mat_Matrix_for_1_for_acc_tmp[2])
          & input_mat_Matrix_for_for_input_mat_Matrix_for_for_nor_3_cse_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1;
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_20_itm_1 <= (input_mat_Matrix_for_1_for_acc_tmp[1])
          & input_mat_Matrix_for_for_input_mat_Matrix_for_for_nor_3_cse_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_rsci_idat <= 17'b00000000000000000;
    end
    else if ( (and_dcpl_89 & exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_4
        & determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_4) | result_rsci_idat_mx0c1
        ) begin
      result_rsci_idat <= MUX_v_17_2_2(determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1,
          determinant_helper_3_do_determinant_ac_int_17_true_determinant_lpi_1, result_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_4
        | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_4) & main_stage_0_5
        ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1 <= determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1 <= 17'b00000000000000000;
    end
    else if ( (mux_nl) & and_dcpl_1 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1 <= nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1[16:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_lpi_1 <= 17'b00000000000000000;
    end
    else if ( main_stage_0_5 & determinant_helper_3_do_determinant_ac_int_17_true_for_and_itm_4
        ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_lpi_1 <= determinant_helper_3_do_determinant_ac_int_17_true_determinant_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_4 <= 1'b0;
    end
    else if ( and_dcpl & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_3_0)
        & exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_3
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_4 <= determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_4
          <= 1'b0;
    end
    else if ( and_dcpl_1 ) begin
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_4
          <= exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_2
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_1_0
          <= 2'b00;
    end
    else if ( and_dcpl_10 ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_2
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_2;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_1_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_3 <=
          1'b0;
    end
    else if ( (mux_3_nl) & main_stage_0_3 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_3 <=
          determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_3
          <= 2'b00;
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_3
          <= 1'b0;
    end
    else if ( and_dcpl_12 ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_3
          <= lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2;
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_3
          <= exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_2
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0
          <= 2'b00;
    end
    else if ( and_dcpl_15 ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_2
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_2;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_2 <=
          1'b0;
    end
    else if ( (mux_5_nl) & main_stage_0_2 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_2 <=
          determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2
          <= 2'b00;
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_2
          <= 1'b0;
    end
    else if ( and_dcpl_17 ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2
          <= lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1;
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_2
          <= exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_2
          <= 1'b0;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0
          <= 2'b00;
    end
    else if ( and_dcpl_20 ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_2
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1;
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0
          <= lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_1_0_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_1 <=
          1'b0;
    end
    else if ( (~((mux_6_nl) | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0))
        | or_dcpl ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_1 <=
          MUX1HOT_s_1_3_2(determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1,
          determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1,
          exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2, {(and_95_nl) , (and_97_nl)
          , or_dcpl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1
          <= 2'b00;
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_1
          <= 1'b0;
    end
    else if ( and_dcpl_22 ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1
          <= lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1;
      exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_1
          <= exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_4;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_Matrix_for_asn_sft_lpi_1 <= 1'b0;
    end
    else if ( ~(input_mat_Matrix_for_for_equal_tmp_2 | input_mat_Matrix_for_for_equal_tmp_3
        | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1)
        ) begin
      input_mat_Matrix_for_asn_sft_lpi_1 <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 <= 1'b0;
    end
    else if ( ~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
        ) begin
      lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 <= lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0 <= 1'b0;
    end
    else if ( ~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
        ) begin
      lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0 <= lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_0_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_Matrix_for_for_j_1_1_1_lpi_1 <= 1'b0;
    end
    else if ( ~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1
        ) begin
      input_mat_Matrix_for_for_j_1_1_1_lpi_1 <= (input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1
          | input_mat_Matrix_for_for_input_mat_Matrix_for_for_nor_3_cse_1) & (lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_1_1
          | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_dfm_3_0_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 <= 1'b0;
    end
    else if ( or_dcpl_4 & (determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1
        | determinant_helper_3_do_determinant_ac_int_17_true_for_and_6_m1c_1) ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 <= MUX_s_1_2_2((input_mat_Matrix_for_input_mat_Matrix_for_and_8_nl),
          (determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_or_nl),
          determinant_helper_3_do_determinant_ac_int_17_true_for_and_6_m1c_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_31_2_lpi_1 <=
          30'b000000000000000000000000000000;
    end
    else if ( (~ (mux_44_nl)) & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
        & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        & nor_85_cse ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_31_2_lpi_1 <=
          MUX_v_30_2_2((determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_and_nl),
          (z_out_3[30:1]), determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_6_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1 <= 1'b0;
    end
    else if ( ~((~((determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1
        & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_or_tmp_1) | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_8_rgt))
        | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
        | or_dcpl_41) ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1 <= MUX_s_1_2_2(determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1,
          (z_out_3[0]), determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_8_rgt);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1 <= 1'b0;
    end
    else if ( ~((~(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4
        | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_13_rgt)) |
        (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
        | or_dcpl_41) ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1 <= MUX_s_1_2_2((determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_9_nl),
          (determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_or_1_nl),
          determinant_helper_3_get_minor_ac_int_17_true_for_and_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1 <= 1'b0;
      determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1 <= 1'b0;
    end
    else if ( determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_and_cse
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1 <= (determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_nl)
          | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3;
      determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1 <= MUX_s_1_2_2((determinant_helper_3_get_minor_ac_int_17_true_for_for_mux_4_nl),
          determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1,
          determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_nor_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
          <= 1'b0;
    end
    else if ( or_dcpl_4 ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
          <= ((determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_2_nl)
          & (~(determinant_helper_3_do_determinant_ac_int_17_true_for_and_25_ssc_1
          | determinant_helper_3_get_minor_ac_int_17_true_for_and_25_ssc_1))) | determinant_helper_3_get_minor_ac_int_17_true_for_and_44_ssc_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0
          <= 2'b00;
    end
    else if ( (~ (mux_10_nl)) | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva
        ) begin
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0
          <= MUX_v_2_2_2((determinant_helper_3_do_determinant_ac_int_17_true_for_and_28_nl),
          2'b11, determinant_helper_3_get_minor_ac_int_17_true_for_and_25_ssc_1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1
          <= 2'b00;
    end
    else if ( ~((mux_46_nl) | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        ) begin
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1
          <= determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1 <= 1'b0;
    end
    else if ( determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
        & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3 & (~
        (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]))
        & (~ or_dcpl_41) ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1 <= determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_dfm_1
          <= 17'b00000000000000000;
    end
    else if ( (determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_4
        | determinant_helper_3_do_determinant_ac_int_17_true_for_or_45_itm_4 | (~
        main_stage_0_5) | determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_3)
        & determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_3 & main_stage_0_4
        ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_dfm_1
          <= MUX_v_17_2_2(17'b00000000000000000, determinant_helper_3_do_determinant_ac_int_17_true_determinant_1_lpi_1_mx0,
          (input_mat_Matrix_for_not_17_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_3
          <= 17'b00000000000000000;
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1
          <= 17'b00000000000000000;
    end
    else if ( and_dcpl_26 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_3
          <= determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1
          <= nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1[16:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      sfi_exit_input_mat_Matrix_for_lpi_1 <= 1'b0;
    end
    else if ( or_dcpl_4 & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_1_1)
        ) begin
      sfi_exit_input_mat_Matrix_for_lpi_1 <= ~((~(sfi_exit_input_mat_Matrix_for_lpi_1
          | input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1)) | input_mat_Matrix_for_for_equal_tmp_2);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_3 <= 1'b0;
    end
    else if ( and_dcpl_9 & exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_2
        & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_3 <= determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_itm_1
          <= 17'b00000000000000000;
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1
          <= 17'b00000000000000000;
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_2
          <= 17'b00000000000000000;
    end
    else if ( and_dcpl_29 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_itm_1
          <= MUX_v_17_2_2((determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_nl),
          determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_1,
          lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[1]);
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1
          <= nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1[16:0];
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_2
          <= MUX_v_17_2_2(determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_1,
          determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_acc_itm_1,
          lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[1]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_2 <= 1'b0;
    end
    else if ( and_dcpl_14 & exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_st_1
        & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_2 <= determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_acc_1_itm_1
          <= 17'b00000000000000000;
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_1
          <= 17'b00000000000000000;
      determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_acc_itm_1
          <= 17'b00000000000000000;
    end
    else if ( and_dcpl_32 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_acc_1_itm_1
          <= nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_ac000000[16:0];
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_1
          <= MUX1HOT_v_17_3_2(input_mat_data_0_2_lpi_1, input_mat_data_0_0_lpi_1,
          (determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_nl),
          {(and_100_nl) , (and_101_nl) , (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]))});
      determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_acc_itm_1
          <= MUX_v_17_2_2((z_out_3[16:0]), determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_0_lpi_1,
          lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1
        | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1) & main_stage_0_2
        & nor_85_cse & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
        & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
        & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0==2'b00)
        & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
        & (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1 <= determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1 <= 17'b00000000000000000;
    end
    else if ( and_dcpl_36 & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0==2'b00)
        & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
        & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
        & nor_85_cse ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_1 <= 1'b0;
    end
    else if ( and_dcpl_36 & or_125_cse & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0==2'b00)
        & determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
        & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
        & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]))
        & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_51_itm_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_1
          & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (~(determinant_helper_3_get_minor_ac_int_17_true_for_or_28_itm_1 &
        determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1))
        & (~ determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1)
        & main_stage_0_2 ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_2_0_lpi_1 <= 17'b00000000000000000;
    end
    else if ( ~((~(and_dcpl_48 | (~ (input_mat_Matrix_for_1_for_acc_tmp[1])))) |
        or_dcpl_42) ) begin
      input_mat_data_2_0_lpi_1 <= input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1
          <= 17'b00000000000000000;
    end
    else if ( or_125_cse & (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
        & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[1])
        & or_dcpl_10 & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1
        & (~ (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[0]))
        & and_dcpl_51 & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31
        & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
        & nor_85_cse ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1
          <= determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_40_itm_1 <= 1'b0;
      determinant_helper_3_get_minor_ac_int_17_true_for_and_41_itm_1 <= 1'b0;
    end
    else if ( determinant_helper_3_get_minor_ac_int_17_true_for_or_33_cse ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_and_40_itm_1 <= MUX_s_1_2_2(determinant_helper_3_get_minor_ac_int_17_true_for_and_36_cse_mx0w0,
          (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]),
          and_dcpl_109);
      determinant_helper_3_get_minor_ac_int_17_true_for_and_41_itm_1 <= MUX_s_1_2_2(determinant_helper_3_get_minor_ac_int_17_true_for_and_28_cse_1,
          (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]),
          and_dcpl_109);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_2_1_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (mux_47_nl) & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        & main_stage_0_2 & determinant_helper_3_do_determinant_ac_int_17_true_for_and_11_itm_1
        ) begin
      input_mat_data_2_1_lpi_1 <= input_mat_data_2_1_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_2_2_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (~(or_177_cse & (input_mat_Matrix_for_1_for_acc_tmp[2]))) & main_stage_0_2
        & determinant_helper_3_do_determinant_ac_int_17_true_for_and_21_itm_1 ) begin
      input_mat_data_2_2_lpi_1 <= input_mat_data_2_2_lpi_1_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1 <= 1'b0;
    end
    else if ( ((~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]))
        | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
        | nand_8_cse | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
        | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
        | nor_11_cse) & or_dcpl_10 & and_dcpl_22 ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1 <= determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_2_itm_1
          <= 17'b00000000000000000;
    end
    else if ( (~ (mux_51_nl)) & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
        & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)
        & (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[0]) ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_2_itm_1
          <= MUX1HOT_v_17_3_2(input_mat_data_1_1_lpi_1, determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_2,
          determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_2_input_mat_getElement_1_slc_input_mat_data_17_16_0_ctmp_sva_1_mx0,
          {(determinant_helper_3_get_minor_ac_int_17_true_for_and_52_nl) , (determinant_helper_3_get_minor_ac_int_17_true_for_or_26_nl)
          , determinant_helper_3_get_minor_ac_int_17_true_for_and_30_cse_1});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1 <= 1'b0;
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1 <= 1'b0;
    end
    else if ( and_dcpl_73 ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1 <= determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
      determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1 <= determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_3;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg
          <= 1'b0;
    end
    else if ( and_dcpl_68 & or_dcpl_10 & input_mat_Matrix_for_i_1_1_lpi_1 & (~ lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1)
        & input_mat_Matrix_for_for_j_1_1_1_lpi_1 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
        ) begin
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_1_dfm_1_reg
          <= ~ exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_dfm_6_1
          <= 17'b00000000000000000;
    end
    else if ( (mux_58_nl) & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
        & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        & (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_dfm_6_1
          <= MUX_v_17_2_2(17'b00000000000000000, (determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_1_nl),
          determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_3);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp <= 1'b0;
    end
    else if ( (((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
        & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
        & (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0==2'b00)
        & determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
        & (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[0])) |
        (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[1])) & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
        & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]))
        & (~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
        | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva))
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp <= determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_4_psp_mx0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_0_lpi_1 <= 17'b00000000000000000;
    end
    else if ( ~((mux_65_nl) | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        ) begin
      determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_0_lpi_1 <= MUX_v_17_2_2(17'b00000000000000000,
          (mux1h_nl), (not_235_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_0_0_lpi_1 <= 17'b00000000000000000;
    end
    else if ( ~(and_dcpl_48 | or_62_cse | (input_mat_Matrix_for_1_for_acc_tmp[0]))
        ) begin
      input_mat_data_0_0_lpi_1 <= input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_0_2_lpi_1 <= 17'b00000000000000000;
    end
    else if ( ~(and_dcpl_48 | or_62_cse | (~ (input_mat_Matrix_for_1_for_acc_tmp[0])))
        ) begin
      input_mat_data_0_2_lpi_1 <= input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1
          <= 17'b00000000000000000;
    end
    else if ( or_177_cse & or_62_cse ) begin
      input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1
          <= input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1
          <= 17'b00000000000000000;
    end
    else if ( (~(or_122_cse & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0))
        & and_dcpl_69 ) begin
      input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1
          <= input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_11_itm_1 <= 1'b0;
    end
    else if ( ~((mux_32_nl) | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        ) begin
      determinant_helper_3_do_determinant_ac_int_17_true_for_and_11_itm_1 <= input_mat_Matrix_for_i_1_1_lpi_1_dfm_1
          & (~ input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1) & (~(input_mat_Matrix_for_for_equal_tmp_2
          | input_mat_Matrix_for_for_equal_tmp_3 | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2
          | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_3));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_1_1_lpi_1 <= 17'b00000000000000000;
      input_mat_data_1_0_lpi_1 <= 17'b00000000000000000;
    end
    else if ( input_mat_data_and_3_cse ) begin
      input_mat_data_1_1_lpi_1 <= input_rsci_idat[84:68];
      input_mat_data_1_0_lpi_1 <= input_rsci_idat[67:51];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_1_2_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (mux_38_nl) & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva)
        & (~(or_dcpl_57 | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)))
        ) begin
      input_mat_data_1_2_lpi_1 <= input_rsci_idat[101:85];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      input_mat_data_0_1_lpi_1 <= 17'b00000000000000000;
    end
    else if ( (~((or_122_cse & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)
        | or_tmp_44)) | exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva
        ) begin
      input_mat_data_0_1_lpi_1 <= input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_exs_34_16_0_ctmp_sva_1_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1_dfm_1_reg
          <= 1'b0;
    end
    else if ( (mux_20_nl) & and_dcpl_69 & (~ lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1)
        & input_mat_Matrix_for_for_j_1_1_1_lpi_1 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
        ) begin
      reg_determinant_helper_3_get_minor_ac_int_17_true_minor_data_1_1_lpi_1_dfm_1_reg
          <= ~ exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2;
    end
  end
  assign input_mat_Matrix_for_for_input_mat_Matrix_for_for_mux_22_nl = MUX_s_1_2_2(input_mat_Matrix_for_i_1_1_lpi_1_dfm_1,
      z_out_1, input_mat_Matrix_for_for_equal_tmp_2);
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_mul_2_itm_1
      = $signed(determinant_helper_3_do_determinant_ac_int_17_true_for_1_input_mat_getElement_2_input_mat_getElement_2_mux_1_itm_3)
      * $signed(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1);
  assign nor_43_nl = ~((~ determinant_helper_3_do_determinant_ac_int_17_true_for_and_12_itm_3)
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_3!=2'b10));
  assign nor_44_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_3[1])
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_1_0[0])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_3_1_0[1]));
  assign mux_nl = MUX_s_1_2_2((nor_43_nl), (nor_44_nl), determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_3);
  assign nor_41_nl = ~((lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0[1])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_2_1_0[0])
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0);
  assign nor_42_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2[0])
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_0);
  assign mux_2_nl = MUX_s_1_2_2((nor_41_nl), (nor_42_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_2[1]);
  assign mux_3_nl = MUX_s_1_2_2(determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_2,
      (mux_2_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_2_1);
  assign nor_39_nl = ~((lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0[1])
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_st_1_1_0[0])
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0);
  assign nor_40_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[0])
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_0);
  assign mux_4_nl = MUX_s_1_2_2((nor_39_nl), (nor_40_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[1]);
  assign mux_5_nl = MUX_s_1_2_2(determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1,
      (mux_4_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_st_1_1);
  assign and_95_nl = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]))
      & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign and_97_nl = and_dcpl_95 & (~ exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_sva);
  assign or_9_nl = (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]));
  assign mux_6_nl = MUX_s_1_2_2((or_9_nl), (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]),
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]);
  assign input_mat_Matrix_for_input_mat_Matrix_for_and_8_nl = determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1
      & (~ exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_or_nl
      = determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_not_4_nl
      = ~ determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_and_nl
      = MUX_v_30_2_2(30'b000000000000000000000000000000, determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_31_2_lpi_1,
      (determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_not_4_nl));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_mux_4_nl = MUX_s_1_2_2((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]),
      determinant_helper_3_get_minor_ac_int_17_true_for_and_41_itm_1, or_dcpl_41);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_6_nl = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4 & (~
      (determinant_helper_3_get_minor_ac_int_17_true_for_mux_4_nl)) & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2;
  assign or_130_nl = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[0])
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31);
  assign and_187_nl = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[1])
      & (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign mux_43_nl = MUX_s_1_2_2(nor_tmp_10, (or_130_nl), and_187_nl);
  assign or_129_nl = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
      | nor_tmp_10;
  assign mux_44_nl = MUX_s_1_2_2((mux_43_nl), (or_129_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_9_nl
      = determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_or_1_nl
      = determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1 | determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_itm_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_nl = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_13_rgt
      & (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]));
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_12_nl = determinant_helper_3_get_minor_ac_int_17_true_for_for_or_3_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_nl = MUX_s_1_2_2(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1,
      determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1, determinant_helper_3_get_minor_ac_int_17_true_for_for_1_and_12_nl);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_or_nl
      = determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_2_acc_itm_2;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_for_mux_4_nl = MUX_s_1_2_2(determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1_dfm_1,
      (determinant_helper_3_get_minor_ac_int_17_true_for_for_determinant_helper_3_get_minor_ac_int_17_true_for_for_or_nl),
      determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_nor_1_nl
      = ~((~(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_4
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5 | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1)) | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | or_dcpl);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_2_nl
      = MUX1HOT_s_1_3_2(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2,
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_dfm_2_1,
      (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1),
      {determinant_helper_3_do_determinant_ac_int_17_true_for_or_47_ssc_1 , determinant_helper_3_do_determinant_ac_int_17_true_for_and_26_ssc_1
      , determinant_helper_3_do_determinant_ac_int_17_true_for_and_27_ssc_1});
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_nor_1_nl = ~(determinant_helper_3_get_minor_ac_int_17_true_for_and_44_ssc_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_and_27_ssc_1);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_28_nl = MUX_v_2_2_2(2'b00,
      determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_1_tmp,
      (determinant_helper_3_do_determinant_ac_int_17_true_for_nor_1_nl));
  assign and_120_nl = ((~ lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1) | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0)
      & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign and_121_nl = input_mat_Matrix_for_for_j_1_1_1_lpi_1 & input_mat_Matrix_for_i_1_1_lpi_1;
  assign mux_8_nl = MUX_s_1_2_2(nor_tmp, (and_120_nl), and_121_nl);
  assign or_17_nl = nor_11_cse | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1!=2'b01)
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0;
  assign mux_9_nl = MUX_s_1_2_2((mux_8_nl), (or_17_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign mux_7_nl = MUX_s_1_2_2(nor_tmp, lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0,
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign or_15_nl = (determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp!=2'b00);
  assign mux_10_nl = MUX_s_1_2_2((mux_9_nl), (mux_7_nl), or_15_nl);
  assign nor_79_nl = ~(nor_11_cse | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | nand_21_cse);
  assign mux_45_nl = MUX_s_1_2_2((nor_79_nl), (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]),
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]);
  assign nand_20_nl = ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1
      & (~ (mux_45_nl)));
  assign or_178_nl = (~ input_mat_Matrix_for_i_1_1_lpi_1) | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1
      | (~ input_mat_Matrix_for_for_j_1_1_1_lpi_1) | lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1;
  assign mux_46_nl = MUX_s_1_2_2((nand_20_nl), (or_178_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign input_mat_Matrix_for_not_17_nl = ~ determinant_helper_3_do_determinant_ac_int_17_true_for_asn_sft_lpi_1_st_3;
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_acc_2_itm_1
      = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_itm_1
      + determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1;
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_nl
      = $signed(determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1)
      * $signed(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_mux_12_itm_1);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_1_nl[16:0];
  assign determinant_helper_2_do_determinant_ac_int_17_true_for_mux_6_nl = MUX_v_17_2_2(determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_acc_itm_1,
      input_mat_data_2_0_lpi_1, lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1_st_1[1]);
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_mul_1_itm_1
      = $signed(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_acc_1_itm_1)
      * $signed(conv_u2s_17_18(determinant_helper_2_do_determinant_ac_int_17_true_for_mux_6_nl));
  assign determinant_helper_2_do_determinant_ac_int_17_true_for_mux_7_nl = MUX_v_17_2_2((~
      input_mat_data_1_2_lpi_1), (~ determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_1_lpi_2),
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_2_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_determinant_helper_2_do_determinant_ac_int_17_true_for_ac000000
      = (determinant_helper_2_do_determinant_ac_int_17_true_for_mux_7_nl) + 17'b00000000000000001;
  assign nl_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_nl
      = $signed(input_mat_data_1_0_lpi_1) * $signed(input_mat_data_2_2_lpi_1_mx0);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_nl
      = nl_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_2_do_determinant_ac_int_17_true_for_1_mul_nl[16:0];
  assign and_100_nl = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
      & determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1;
  assign and_101_nl = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0])
      & (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1);
  assign nor_73_nl = ~((~ input_mat_Matrix_for_i_1_1_lpi_1) | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1
      | (~(input_mat_Matrix_for_for_j_1_1_1_lpi_1 & lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)));
  assign nor_74_nl = ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
      | (~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | nor_11_cse | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | nand_21_cse)));
  assign mux_47_nl = MUX_s_1_2_2((nor_73_nl), (nor_74_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_52_nl = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1)
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_26_nl = (determinant_helper_3_get_minor_ac_int_17_true_for_for_or_2_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1) | determinant_helper_3_get_minor_ac_int_17_true_for_and_29_cse_1
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_5 | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1 | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]);
  assign or_153_nl = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | not_tmp_119;
  assign and_184_nl = (determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[0]))
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1 & determinant_helper_3_get_minor_ac_int_17_true_for_unequal_tmp_1_1;
  assign mux_48_nl = MUX_s_1_2_2(not_tmp_119, (and_184_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[1]);
  assign or_150_nl = (~((lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1))) |
      nor_tmp_15;
  assign mux_49_nl = MUX_s_1_2_2((mux_48_nl), (or_150_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2);
  assign mux_50_nl = MUX_s_1_2_2((mux_49_nl), nor_tmp_15, lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]);
  assign mux_51_nl = MUX_s_1_2_2((or_153_nl), (mux_50_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_45_nl = (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_or_tmp_1)
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_or_25_nl = (determinant_helper_3_get_minor_ac_int_17_true_for_for_or_tmp_1
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1) | determinant_helper_3_get_minor_ac_int_17_true_for_and_29_cse_1
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_equal_tmp_3 | determinant_helper_3_get_minor_ac_int_17_true_for_for_1_nor_tmp_1
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | ((~ and_182_cse) & determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_48_nl = and_182_cse
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_11_m1c_1;
  assign determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_1_nl
      = MUX1HOT_v_17_4_2(input_mat_data_1_0_lpi_1, determinant_helper_3_get_minor_ac_int_17_true_minor_data_0_0_lpi_1_mx0,
      input_mat_data_1_1_lpi_1, input_mat_data_2_2_lpi_1_mx0, {(determinant_helper_3_get_minor_ac_int_17_true_for_and_45_nl)
      , (determinant_helper_3_get_minor_ac_int_17_true_for_or_25_nl) , determinant_helper_3_get_minor_ac_int_17_true_for_and_30_cse_1
      , (determinant_helper_3_get_minor_ac_int_17_true_for_and_48_nl)});
  assign nand_13_nl = ~(((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1!=2'b10))
      & (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[1]));
  assign or_161_nl = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2
      | (~ main_stage_0_2) | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  assign or_160_nl = (~(determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_1_lpi_1
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2)))
      | (~ main_stage_0_2) | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  assign or_159_nl = (~(determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1
      | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31)))
      | (~ main_stage_0_2) | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  assign or_158_nl = and_182_cse | (~ main_stage_0_2) | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  assign mux_53_nl = MUX_s_1_2_2((or_159_nl), (or_158_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[0]);
  assign mux_54_nl = MUX_s_1_2_2((or_160_nl), (mux_53_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[1]);
  assign and_183_nl = nand_8_cse & or_tmp_77;
  assign or_155_nl = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00);
  assign mux_52_nl = MUX_s_1_2_2((and_183_nl), or_tmp_77, or_155_nl);
  assign mux_55_nl = MUX_s_1_2_2((mux_54_nl), (mux_52_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2);
  assign mux_56_nl = MUX_s_1_2_2((or_161_nl), (mux_55_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign or_154_nl = (~ (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]))
      | (~ main_stage_0_2) | determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_1_1
      | determinant_helper_3_do_determinant_ac_int_17_true_for_or_tmp_1_1;
  assign mux_57_nl = MUX_s_1_2_2((mux_56_nl), (or_154_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1]);
  assign mux_58_nl = MUX_s_1_2_2((nand_13_nl), (mux_57_nl), determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[0]);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_33_nl = determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2
      & determinant_helper_3_get_minor_ac_int_17_true_for_and_9_m1c_1 & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2
      & (~ and_128_tmp);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_56_nl = (~ or_dcpl_42)
      & determinant_helper_3_get_minor_ac_int_17_true_for_or_32_m1c & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2
      & (~ and_128_tmp);
  assign determinant_helper_3_get_minor_ac_int_17_true_for_and_57_nl = or_dcpl_42
      & determinant_helper_3_get_minor_ac_int_17_true_for_or_32_m1c & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2
      & (~ and_128_tmp);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_and_35_nl = determinant_helper_3_get_minor_ac_int_17_true_for_and_28_cse_1
      & determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2 & (~ and_128_tmp);
  assign mux1h_nl = MUX1HOT_v_17_5_2((signext_17_1(~ exit_input_mat_Matrix_for_lpi_1_dfm_3_mx0w2)),
      input_mat_data_1_2_lpi_1, input_mat_Matrix_for_for_slc_input_mat_Matrix_for_for_acc_psp_1_34_16_0_ctmp_sva_1,
      input_mat_data_2_0_lpi_1, input_mat_data_2_1_lpi_1_mx0, {(~ determinant_helper_3_do_determinant_ac_int_17_true_for_equal_tmp_2)
      , (determinant_helper_3_get_minor_ac_int_17_true_for_and_33_nl) , (determinant_helper_3_get_minor_ac_int_17_true_for_and_56_nl)
      , (determinant_helper_3_get_minor_ac_int_17_true_for_and_57_nl) , (determinant_helper_3_do_determinant_ac_int_17_true_for_and_35_nl)});
  assign not_235_nl = ~ and_128_tmp;
  assign or_179_nl = (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0)
      | lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_1 | (~(input_mat_Matrix_for_for_j_1_1_1_lpi_1
      & input_mat_Matrix_for_i_1_1_lpi_1));
  assign nor_82_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | (~ (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[1])));
  assign mux_63_nl = MUX_s_1_2_2((nor_82_nl), (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[1]),
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign nor_83_nl = ~((lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2);
  assign or_168_nl = determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[0]);
  assign mux_60_nl = MUX_s_1_2_2((~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_acc_itm_2),
      (or_168_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2);
  assign nand_23_nl = ~(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_1_for_1_1_acc_itm_31
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1);
  assign or_166_nl = (~ determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_1_acc_itm_2)
      | determinant_helper_3_get_minor_ac_int_17_true_for_for_col_1_lpi_1 | (~(determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_acc_itm_2
      | determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1 | (determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[1])));
  assign mux_59_nl = MUX_s_1_2_2((nand_23_nl), (or_166_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[0]);
  assign or_167_nl = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
      | (mux_59_nl);
  assign mux_61_nl = MUX_s_1_2_2((mux_60_nl), (or_167_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0[1]);
  assign or_169_nl = (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[1])
      | (mux_61_nl);
  assign mux_62_nl = MUX_s_1_2_2((nor_83_nl), (or_169_nl), lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign mux_64_nl = MUX_s_1_2_2((mux_63_nl), (mux_62_nl), determinant_helper_3_get_minor_ac_int_17_true_for_mux1h_24_tmp[0]);
  assign or_180_nl = lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
      | (mux_64_nl);
  assign mux_65_nl = MUX_s_1_2_2((or_179_nl), (or_180_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign mux_32_nl = MUX_s_1_2_2((~ mux_31_itm), or_tmp_41, lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0);
  assign mux_36_nl = MUX_s_1_2_2(sfi_exit_input_mat_Matrix_for_lpi_1, (~ input_mat_Matrix_for_i_1_1_lpi_1),
      input_mat_Matrix_for_asn_sft_lpi_1);
  assign nor_15_nl = ~(lfst_exitL_exit_input_mat_Matrix_for_2_for_lpi_1_0 | (mux_36_nl));
  assign mux_37_nl = MUX_s_1_2_2(input_mat_Matrix_for_i_1_1_lpi_1, (nor_15_nl), and_124_cse);
  assign nor_16_nl = ~(lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_0
      | (~(nor_11_cse | (~ determinant_helper_3_do_determinant_ac_int_17_true_for_j_1_lpi_1)
      | (~ determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1)
      | (lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1!=2'b01)
      | (~ lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2)
      | (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_1_0!=2'b00))));
  assign mux_38_nl = MUX_s_1_2_2((mux_37_nl), (nor_16_nl), lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_lpi_1_dfm_3_1);
  assign nor_23_nl = ~((determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp[1])
      | (~ and_dcpl_51));
  assign mux_18_nl = MUX_s_1_2_2(and_dcpl_51, determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1,
      lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2);
  assign or_47_nl = (lfst_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_1_determinant_helper_3_get_minor_ac_int_17_true_for_2_for_2_lpi_1_2
      & determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_5_1_lpi_1) |
      and_dcpl_51;
  assign or_46_nl = (determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp[1])
      | (determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_1_tmp!=2'b00);
  assign mux_19_nl = MUX_s_1_2_2((mux_18_nl), (or_47_nl), or_46_nl);
  assign mux_20_nl = MUX_s_1_2_2((nor_23_nl), (mux_19_nl), determinant_helper_3_do_determinant_ac_int_17_true_for_mux1h_42_tmp[0]);
  assign determinant_helper_3_do_determinant_ac_int_17_true_for_mux_15_nl = MUX_v_31_2_2((signext_31_17(~
      input_mat_data_0_1_lpi_1)), ({determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_31_2_lpi_1
      , determinant_helper_3_get_minor_ac_int_17_true_for_for_1_col2_7_1_lpi_1}),
      lfst_exitL_exit_determinant_helper_3_do_determinant_ac_int_17_true_for_2_determinant_helper_3_get_minor_ac_int_17_true_for_lpi_1[0]);
  assign nl_z_out_3 = (determinant_helper_3_do_determinant_ac_int_17_true_for_mux_15_nl)
      + 31'b0000000000000000000000000000001;
  assign z_out_3 = nl_z_out_3[30:0];
  assign input_mat_Matrix_for_for_input_mat_Matrix_for_for_or_6_nl = input_mat_Matrix_for_i_1_1_lpi_1_dfm_1
      | (~ sfi_exit_input_mat_Matrix_for_lpi_1);
  assign input_mat_Matrix_for_for_mux_25_nl = MUX_s_1_2_2(input_mat_Matrix_for_asn_sft_lpi_1,
      (input_mat_Matrix_for_for_input_mat_Matrix_for_for_or_6_nl), and_dcpl_121);
  assign input_mat_Matrix_for_for_mux_26_nl = MUX_s_1_2_2(input_mat_Matrix_for_for_j_1_1_1_lpi_1_dfm_1,
      input_mat_Matrix_for_asn_sft_lpi_1, and_dcpl_121);
  assign z_out_1 = MUX_s_1_2_2((input_mat_Matrix_for_for_mux_25_nl), input_mat_Matrix_for_i_1_1_lpi_1_dfm_1,
      input_mat_Matrix_for_for_mux_26_nl);

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_3_2;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [2:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    MUX1HOT_v_17_3_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_4_2;
    input [16:0] input_3;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [3:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    result = result | ( input_3 & {17{sel[3]}});
    MUX1HOT_v_17_4_2 = result;
  end
  endfunction


  function automatic [16:0] MUX1HOT_v_17_5_2;
    input [16:0] input_4;
    input [16:0] input_3;
    input [16:0] input_2;
    input [16:0] input_1;
    input [16:0] input_0;
    input [4:0] sel;
    reg [16:0] result;
  begin
    result = input_0 & {17{sel[0]}};
    result = result | ( input_1 & {17{sel[1]}});
    result = result | ( input_2 & {17{sel[2]}});
    result = result | ( input_3 & {17{sel[3]}});
    result = result | ( input_4 & {17{sel[4]}});
    MUX1HOT_v_17_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | ( input_1 & {2{sel[1]}});
    result = result | ( input_2 & {2{sel[2]}});
    result = result | ( input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_2_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [0:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_17_2_2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_4_2x1x2;
    input [16:0] input_0;
    input [16:0] input_3;
    input [1:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      default : begin
        result = input_3;
      end
    endcase
    MUX_v_17_4_2x1x2 = result;
  end
  endfunction


  function automatic [16:0] MUX_v_17_5_2;
    input [16:0] input_0;
    input [16:0] input_1;
    input [16:0] input_2;
    input [16:0] input_3;
    input [16:0] input_4;
    input [2:0] sel;
    reg [16:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      default : begin
        result = input_4;
      end
    endcase
    MUX_v_17_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [29:0] MUX_v_30_2_2;
    input [29:0] input_0;
    input [29:0] input_1;
    input [0:0] sel;
    reg [29:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_30_2_2 = result;
  end
  endfunction


  function automatic [30:0] MUX_v_31_2_2;
    input [30:0] input_0;
    input [30:0] input_1;
    input [0:0] sel;
    reg [30:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_31_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_32_1_31;
    input [31:0] vector;
    reg [31:0] tmp;
  begin
    tmp = vector >> 31;
    readslicef_32_1_31 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [16:0] signext_17_1;
    input [0:0] vector;
  begin
    signext_17_1= {{16{vector[0]}}, vector};
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [30:0] signext_31_17;
    input [16:0] vector;
  begin
    signext_31_17= {{14{vector[16]}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2s_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2s_2_3 =  {1'b0, vector};
  end
  endfunction


  function automatic [17:0] conv_u2s_17_18 ;
    input [16:0]  vector ;
  begin
    conv_u2s_17_18 =  {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    determinant
// ------------------------------------------------------------------


module determinant (
  clk, rst, input_rsc_dat, input_rsc_triosy_lz, result_rsc_dat, result_rsc_triosy_lz
);
  input clk;
  input rst;
  input [152:0] input_rsc_dat;
  output input_rsc_triosy_lz;
  output [16:0] result_rsc_dat;
  output result_rsc_triosy_lz;



  // Interconnect Declarations for Component Instantiations 
  determinant_core determinant_core_inst (
      .clk(clk),
      .rst(rst),
      .input_rsc_dat(input_rsc_dat),
      .input_rsc_triosy_lz(input_rsc_triosy_lz),
      .result_rsc_dat(result_rsc_dat),
      .result_rsc_triosy_lz(result_rsc_triosy_lz)
    );
endmodule



